magic
tech sky130A
magscale 1 2
timestamp 1677477959
<< error_s >>
rect 864 1680 1040 1708
rect 836 1652 858 1680
rect 856 1552 858 1558
rect 1044 1530 1068 1648
rect 856 1524 886 1530
rect 159 880 261 896
rect 351 880 453 896
rect 858 884 1016 908
rect 187 852 233 868
rect 283 846 329 862
rect 379 852 425 868
rect 255 818 357 834
<< metal1 >>
rect 168 2456 368 2540
rect 8 2264 500 2456
rect 8 2208 792 2264
rect 8 2108 500 2208
rect -228 1992 288 2036
rect -228 1504 -184 1992
rect 622 1888 792 2208
rect 96 1802 792 1888
rect 864 1680 1040 1682
rect 194 1552 858 1680
rect 728 1530 856 1552
rect 1040 1530 1044 1648
rect -480 1426 -280 1504
rect -230 1460 382 1504
rect -228 1426 -184 1460
rect -480 1382 -184 1426
rect -480 1304 -280 1382
rect -228 1048 -184 1382
rect 728 1330 1046 1530
rect -228 1004 286 1048
rect -228 710 -184 1004
rect 728 946 856 1330
rect 104 884 858 946
rect 104 880 1016 884
rect 728 866 856 880
rect 194 770 830 834
rect -228 666 400 710
rect -8 452 492 614
rect 654 452 820 770
rect -8 388 824 452
rect -8 348 492 388
rect 220 244 420 348
use sky130_fd_pr__nfet_01v8_H3H3JC  XM1
timestamp 1677474599
transform 1 0 258 0 1 857
box -311 -310 311 310
use sky130_fd_pr__pfet_01v8_3YVXDD  XM2
timestamp 1677474599
transform 1 0 257 0 1 1755
box -311 -419 311 419
<< labels >>
flabel metal1 -480 1304 -280 1504 0 FreeSans 256 0 0 0 in
port 0 nsew
flabel metal1 846 1330 1046 1530 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 168 2340 368 2540 0 FreeSans 256 0 0 0 vdd
port 2 nsew
flabel metal1 220 244 420 444 0 FreeSans 256 0 0 0 vss
port 3 nsew
<< end >>
