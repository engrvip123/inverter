** sch_path: /home/vipul/inverter/xschem/inverter_tb.sch
**.subckt inverter_tb out
*.opin out
x1 vdd inp out GND inverter
VDD vdd GND 1.8
Vinp inp GND PWL(0 0 200n 0 300n 1.8 500n 1.8 600n 0)
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.control
tran 1n 1u
plot V(inp) V(out)
.endc

**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/vipul/inverter/xschem/inverter.sym
** sch_path: /home/vipul/inverter/xschem/inverter.sch
.subckt inverter  vdd in out vss
*.ipin in
*.opin out
*.ipin vdd
*.ipin vss
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.4 W=4 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.4 W=4 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
