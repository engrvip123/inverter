magic
tech sky130A
magscale 1 2
timestamp 1677474599
<< error_p >>
rect -29 172 29 178
rect -29 138 -17 172
rect -29 132 29 138
rect -125 -138 -67 -132
rect 67 -138 125 -132
rect -125 -172 -113 -138
rect 67 -172 79 -138
rect -125 -178 -67 -172
rect 67 -178 125 -172
<< pwell >>
rect -311 -310 311 310
<< nmos >>
rect -111 -100 -81 100
rect -15 -100 15 100
rect 81 -100 111 100
<< ndiff >>
rect -173 88 -111 100
rect -173 -88 -161 88
rect -127 -88 -111 88
rect -173 -100 -111 -88
rect -81 88 -15 100
rect -81 -88 -65 88
rect -31 -88 -15 88
rect -81 -100 -15 -88
rect 15 88 81 100
rect 15 -88 31 88
rect 65 -88 81 88
rect 15 -100 81 -88
rect 111 88 173 100
rect 111 -88 127 88
rect 161 -88 173 88
rect 111 -100 173 -88
<< ndiffc >>
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
<< psubdiff >>
rect -275 240 -179 274
rect 179 240 275 274
rect -275 178 -241 240
rect 241 178 275 240
rect -275 -240 -241 -178
rect 241 -240 275 -178
rect -275 -274 -179 -240
rect 179 -274 275 -240
<< psubdiffcont >>
rect -179 240 179 274
rect -275 -178 -241 178
rect 241 -178 275 178
rect -179 -274 179 -240
<< poly >>
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -111 100 -81 126
rect -33 122 33 138
rect -15 100 15 122
rect 81 100 111 126
rect -111 -122 -81 -100
rect -129 -138 -63 -122
rect -15 -126 15 -100
rect 81 -122 111 -100
rect -129 -172 -113 -138
rect -79 -172 -63 -138
rect -129 -188 -63 -172
rect 63 -138 129 -122
rect 63 -172 79 -138
rect 113 -172 129 -138
rect 63 -188 129 -172
<< polycont >>
rect -17 138 17 172
rect -113 -172 -79 -138
rect 79 -172 113 -138
<< locali >>
rect -275 240 -179 274
rect 179 240 275 274
rect -275 178 -241 240
rect 241 178 275 240
rect -33 138 -17 172
rect 17 138 33 172
rect -161 88 -127 104
rect -161 -104 -127 -88
rect -65 88 -31 104
rect -65 -104 -31 -88
rect 31 88 65 104
rect 31 -104 65 -88
rect 127 88 161 104
rect 127 -104 161 -88
rect -129 -172 -113 -138
rect -79 -172 -63 -138
rect 63 -172 79 -138
rect 113 -172 129 -138
rect -275 -274 -241 -178
rect 241 -274 275 -178
<< viali >>
rect -17 138 17 172
rect -161 1 -127 71
rect -65 -35 -31 35
rect 31 1 65 71
rect 127 -35 161 35
rect -113 -172 -79 -138
rect 79 -172 113 -138
rect -241 -274 -179 -240
rect -179 -274 179 -240
rect 179 -274 241 -240
<< metal1 >>
rect -29 172 29 178
rect -29 138 -17 172
rect 17 138 29 172
rect -29 132 29 138
rect -167 71 -121 83
rect -167 1 -161 71
rect -127 1 -121 71
rect 25 71 71 83
rect -167 -11 -121 1
rect -71 35 -25 47
rect -71 -35 -65 35
rect -31 -35 -25 35
rect 25 1 31 71
rect 65 1 71 71
rect 25 -11 71 1
rect 121 35 167 47
rect -71 -47 -25 -35
rect 121 -35 127 35
rect 161 -35 167 35
rect 121 -47 167 -35
rect -125 -138 -67 -132
rect -125 -172 -113 -138
rect -79 -172 -67 -138
rect -125 -178 -67 -172
rect 67 -138 125 -132
rect 67 -172 79 -138
rect 113 -172 125 -138
rect 67 -178 125 -172
rect -253 -240 253 -234
rect -253 -274 -241 -240
rect 241 -274 253 -240
rect -253 -280 253 -274
<< properties >>
string FIXED_BBOX -258 -257 258 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 40 viadrn -40 viagate 100 viagb 100 viagr 0 viagl 0 viagt 0
<< end >>
